///////////////////////////////////////////////////////////////////////////////////
// Filename:ddr_assertion.sv
// 
// Author: Scaledge
// Date: 24/12/2025
// Revision: 1
// Company: Scaledge Technology Pvt.
// Copyright (c) 2025 Scaledge Technology Pvt. All rights reserved.
// This file is part of the  DDR project.
// Description:
// Dependencies:
// Notes:
//////////////////////////////////////////////////////////////////////////

`ifndef DDR_ASSERTION_SV
`define DDR_ASSERTION_SV

module ddr_assertion(ddr_interface inf);

endmodule

`endif
