///////////////////////////////////////////////////////////////////////////////////
// Filename:ddr_defines.sv
// 
// Author: Scaledge
// Date: 24/12/2025
// Revision: 1
// 
// Company: Scaledge Technology Pvt.
// 
// Copyright (c) <Year> Scaledge Technology Pvt. All rights reserved.
// 
// This file is part of the  VIP project.
// Description:
// Dependencies:
// Notes:
//////////////////////////////////////////////////////////////////////////////////

`define TIMEPERIOD 2.5 //((1/(FREQUENCY))*(1000)) = (1/400)*1000 frq in MHZ 
`define MEM_DQ_WIDTH 8
`define MEM_BA_WIDTH 3
`define MEM_ROW_WIDTH 13
`define MEM_COL_WIDTH 13
`define AL 3
`define CWL 5
`define CL 5
